� �  @                                                                                                                                                                                                                                                 UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUU  UUUUUUUUUUUUUUUU@                                                       UUU  UUUUUUUUUUUUUUUU@                                                       UUU  UUUUUUUUUUUUUUUU@                                                       UUU @UUUUUUUUUUUUUUU@                                                       UUU @UUUUUUUUUUUUUUU@                                                       UUU @UUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                       UUUUUUUUUUUUUUUUUUUUUUU@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      