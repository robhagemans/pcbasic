� �  @                                                                                <     <<���� |                                                                 f      fffbb� �                                                                 0x�8�v 0�fhh� �                                                                 �f� �|xx� |                                                                 |�f| �lhh� �                                                                 f�lf fffbb� �                                                                 <v8<f� <<���� |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       