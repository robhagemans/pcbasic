� �  �>                                                                                                                                                                                                                                                |     8 �     |<���� |                                                       �     l `     �ffff� �                                                       �      l `      ��fbb� �                                                       `x�8�v 8 `|x<8�v `�fhh� �                                                       8�f� v `�lf� 8�|xx� ~                                                       |�f� � `�|�f� �lhh�                                                        ��lf� � b���f� ��fbb�                                                        ��8f� � f���f� �ffff�                                                        |v<f| v �|vv<f| |<���� x                                                                                                                                          x         x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        