� �  @                                                                                 <     8 �     <<���� |                                                       f      l `      fffbb� �                                                       0x�8�v 8 `|x|8�v 0�fhh� �                                                       �f� v `��f� �|xx� |                                                       |�f| � b�|�f| �lhh� �                                                       f�lf � f���f fffbb� �                                                       <v8<f� v �|vv<f� <<���� |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      