� �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                        �                                                                         �     �   0                                                                     0     �   �                                                                     0     �   �                                                                          �   �     0                                                                   �        �                                                                   �                                                                  �         �                                                                  0     �   �  �    0                                                              �   �  �    �     �                                               �         �0   �  2                                                               0   �0   �  2         0                                                 �            ��  8                                                                      ��  �    �                                                       �    �     ��  �        �                                                       0   �  ��         �      �                                             �       ��  ��          8      <                                             �    �   0  �� �   �                                                 �      �   0   0  �� �      2      �                                        �     �0         �        �     <                                                       �                                                               0   ��    � 8   �   �     �                                             0        0  �   � 8     �    <�                                              �     0     �  � �     8                                                 �       ��  0  � �     �    �                                              �     0   0 0  � �  �      >�                                              
 <        ��    �          ?                                   �       �    0  �  � ��       �      <                                      �      (�   �   � � �     �   >      <�                                       <          0 0 # �  � �  �     <�                                               �<   �  � ��   8   �     �                                         ( �    ��  0  ���8  �  >     �                                           
� �    ��  � 00�8     �    �                                               � ?    
  0 � ��  � �  �   �          �                                     
��     � # ���   :   �         �                                         � �   (0 0�#��   �  �        �                                ?�          
�<    � # �À � �  �       ?�*�                                   ��         ��  ���#�� �8 8  �      ?ª                                         ��       
�  � ,��� �� �     ?ʨ                                        �   �      �� ����� � :�    ��                                             ��  �     *? 
�,,"� �8 :    ���                                                   *�� ?�   ��
��.Ȃ *   ��                                                          �� ��  *�+�� �� ��                                                               �����,��(��             ������                                                  
��*����     ?����������                                      
��������������������������                                                 �������                 �����
��                                                                     *� *���
� 
��                                                               ��  +�+��( �   ��                                                          *��   � � �� �� *�     ���                                                   
��    � ,,� � 
�       ���                                              ���     
�   , �����  �         *��                                        *��       +� � ����  
�  *�          *���                                 ��        �   � , ��  � +   �              �                               ��        �   , ���,�  �    ��                                         �          
�   � ,     � �  �    
�                                      �           *�   � � �   ,   �    ��                                                ��    �      �  �  
�     (�                                             ��    +   � , ,   � �    +      
�                                           �     
�    �     � ,  �   �       ��                                        
<     �   � � �   ,       �       (?                                      (�      �       �     �      0        �                                    �      +�   �  , � ,   ,  �   
�         �                                 �      
�      �   , �    ,    +�                                         �      �    ,  �   , � 0  �    �                                                �    �      ,  �  �   ,     �                                               (�    ,      ,  ,  ,     �    <                                             
0    �  �     ,  ,  �   ,     
0                                           �     ,      �  ,     �   �      �                                          �    0   ,   �  ,     #    ,      �                                         �     #    �  �  ,  �  �   �                                              <      �   �  �  ,   �   �    ,                                                             ,   �   #    �                                             �      �    ,   #   ,   ,   �    ,                                            0      �    �   ,      #   0     0                                                      �   �          #                                                       �    #    �      �   �     0                                                     �   0      0   0                                                     �    0   �       �    �      0                                                   �   �       �     �                                                   0                 #     0                                                         0    #                                                                       �             �     �                                                                      �     0                                                             0         0                                                             0     0     �                                                                  �     �     �                                                                        �     �                                                                             �     �                                                                        �                                                                               �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �   0                                                                     �     �   0                                                                     0     �   �                                                                     0     �   �     0                                                         0          �        �                                                                   �                                                                           �                                                                  �     �   �       0                                                                �   �  �    �     0                                                         0   �                                                           0      �   �0   �  2                                                               0       ��  8    8     �                                                 0    �       ��  �    �                                                                 ��  �   �    0                                                   0    0     ��  �                                                               �   ��  ��     8    2                                                    0       ��  �� �   �    �      �                                                 �   0  �� �  �   �     <                                              0   �0    ��        �                                               0               �    8   �     �                                           �    ��   �    � 2   �   2     <�                                           �       �0  �   � 8  �                                                          ��    ��  � 8          �                                              <         �  � �  8   �    >�       �                                      ( �    ��  �� 0  � �  �  �           �                                         �     0 0  �� �  8    �       �                                  �       �    ��   ��   �   >�     �                                    ?      �   
  �� � �� 8  8   �     �                                      �     �0    � 0 # �  �  �   �     �                                        �     
 �     �� �    >     �                                           �         � � ��   �  �    (                                          �      (   �0�8 8    �    �                                             * �     <   �00�  � 8  >    ?�          �                                   � �    ��  � ����� �   >�         �                                       * ?   �� (��,��   �   >�        �                              �          ��  �  �0#��8 � :   ��       ?�*                                 �          *�  
<  �À� �  �       ?���                                     �        �<  
0 ����  �  �      ?¨                                           ?�       �  (���� 8 �     ?ʠ                                          ��   ��     
�� # �,��88 �    �*�                                                
�� ��    �� �.�����   ��                                                       *� �   
� ��Ȼ�8�  ��                                                             ���  �²+����                 ���                                             ���
�ꪊ��        ���������                                                      *�������������                                                ��������������    *����                                                                        
������� ��                                                                   �� ��"� �*   *��                                                            
��  
�(,����
�    *��                                                      ��    *�
 �� 
  �      
��                                                 *��     � � ���+  *�       
���                                          ���     �  � �  ���, �  �         ���                                     ���       
�  +  ��� ,� �   ��            ?�                                �?�        
�  
� � ��  , �   
�                                           �          +�  �  ,   �� 
�   �                                        �           ��   �  � �   , ,  +     +�                                                 �       �    �  �     
�                                               
<    �     ,   �� ,   �     ��                                            (�     �  � , ,   �   �  �      *�                                          ��     /   ,  � �       (   
�      
��                                      ��     �  �   �   , �  �   +�        �                                    �      0   ,   �     �      �         ?                                   ?       �   �  � � ,   #   �    �         �                                <       #      �   , � �      <                                         �       �    �      ,  �  �   �    
�                                       �       <       ,  ,  ,  �  ,        (�                                              �     �   �  ,  ,  ,  �   �     ��                                            #�       �  �  ,     �         �                                           0     �      �  ,     ,    �                                                     �   ,  �  ,  �  �          <                                              �   0  �  ,  �  0    �       �                                       �     �   �     ,   �   �            �                                     <      ,    ,      ,   ,   �    �                                                  0    �   ,      ,   0    �                                                  #    �   ,          �                                                       0        �      �   #      �                                                     ,    �      �   0                                                     0     �   �       �    �      �                                               �    �   �       �    #                                                             �       ,     0                                                    �                 #                                                               0    #                                                                       �             �     �                                                                      0                                                                  0     �    0                                                             0     0     �                                                                        �     �                                                                        �     �                                                                             �     �                                                                         �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     