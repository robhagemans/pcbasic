� �  �>                                                                                                                                                                                                                                                |     |<���� |                                                                 �     �ffff� �                                                                 �      ��fbb� �                                                                 `x�8�v `�fhh� �                                                                 8�f� 8�|xx� ~                                                                 |�f� �lhh�                                                                  ��lf� ��fbb�                                                                  ��8f� �ffff�                                                                  |v<f| |<���� x                                                                                                                                                     x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        