� �  �                                        <     <<���� �                         f      fffbb� �                         0x�8�v 0�fhh�                          �f� �|xx�                          |�f| �lhh� 0                         f�lf fffbb� 0                         <v8<f� <<���� 0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       